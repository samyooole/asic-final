parameter CLK_PERIOD = 10;        // Change based on timing violations from sdf backannotation
parameter PIPE_STAGES = 1;       // Change based on how long it takes to get first output

