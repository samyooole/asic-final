/home/sh2663/asap7_rundir/asic-final/apr/asap7_tech_4x_170803.lef