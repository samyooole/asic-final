/home/sh2663/asap7_rundir/asic-final/apr/asap7sc7p5t_24_R_4x_170912.lef